//=======================================================
//  Title: Lghtweight cosine transform in GF(256) Defines
//=======================================================

`ifndef FF256_LIGHTWEIGHT_COS_TRANSF_DEFINES_V
`define FF256_LIGHTWEIGHT_COS_TRANSF_DEFINES_V

    // FSM defines
    `define IDLE    4'b0000
    `define S0      4'b0001
    `define S1      4'b0010
    `define S2      4'b0011
    `define S3      4'b0100
    `define S4      4'b0101
    `define S5      4'b0110
    `define S6      4'b0111
    `define S7      4'b1000
    `define DONE    4'b1001

`endif