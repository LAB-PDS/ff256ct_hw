//=======================================================
//  Title: Multiplier GF(256) Defines
//=======================================================

`ifndef FF256_LIGHTWEIGHT_COS_TRANSF_DEFINES_V
`define FF256_LIGHTWEIGHT_COS_TRANSF_DEFINES_V

`endif