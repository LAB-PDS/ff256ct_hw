//=======================================================
//  Title: AVALON TO WISHBONE BRIDGE DEFINES
//  Description: Defines used for Avalon/Wishbone interfaces
//=======================================================

`ifndef CUSTOM_RAM_V
`define CUSTOM_RAM_V

// Avalon Memory Mepped Defines
`define AVMM_DATA_WIDTH 32 // Avalon Memory Mapped Data Width
`define AVMM_ADDR_WIDTH 4  // Avalon Memory Mapped Address Width
`define AVMM_BE_WIDTH   4  // Avalon Memory Mapped Byte Enable Width

`endif